`ifndef INSTRUCTION_INCLUDED
`define INSTRUCTION_INCLUDED

typedef enum logic [31:0]{
    SYSCALL = 32'b000000_????????????????????_001100,
    NOP     = 32'b000000_00000000000000000000_000000,
    
    ADD     = 32'b000000_????????????????????_100000,
    ADDU    = 32'b000000_????????????????????_100001,
    SUB     = 32'b000000_????????????????????_100010,
    SUBU    = 32'b000000_????????????????????_100011,
    SLL     = 32'b000000_00000???????????????_000000,
    SRL     = 32'b000000_????????????????????_000010,
    SRA     = 32'b000000_????????????????????_000011,
    SLLV    = 32'b000000_????????????????????_000100,
    SRLV    = 32'b000000_????????????????????_000110,
    SRAV    = 32'b000000_????????????????????_000111,
    AND     = 32'b000000_????????????????????_100100,
    OR      = 32'b000000_????????????????????_100101,
    XOR     = 32'b000000_????????????????????_100110,
    NOR     = 32'b000000_????????????????????_100111,
    SLT     = 32'b000000_????????????????????_101010,
    SLTU    = 32'b000000_????????????????????_101011,

    ADDI    = 32'b001000_????????????????????_??????,
    ADDIU   = 32'b001001_????????????????????_??????,
    ANDI    = 32'b001100_????????????????????_??????,
    ORI     = 32'b001101_????????????????????_??????,
    XORI    = 32'b001110_????????????????????_??????,
    SLTI    = 32'b001010_????????????????????_??????,
    SLTIU   = 32'b001011_????????????????????_??????,

    LUI     = 32'b001111_????????????????????_??????,

    MULT    = 32'b000000_????????????????????_011000,
    MULTU   = 32'b000000_????????????????????_011001,
    DIV     = 32'b000000_????????????????????_011010,
    DIVU    = 32'b000000_????????????????????_011011,
    MFHI    = 32'b000000_????????????????????_010000,
    MTHI    = 32'b000000_????????????????????_010001,
    MFLO    = 32'b000000_????????????????????_010010,
    MTLO    = 32'b000000_????????????????????_010011,

    BEQ     = 32'b000100_????????????????????_??????,
    BNE     = 32'b000101_????????????????????_??????,
    BLEZ    = 32'b000110_????????????????????_??????,
    BGTZ    = 32'b000111_????????????????????_??????,
    BGEZ    = 32'b000001_?????00001??????????_??????,
    BLTZ    = 32'b000001_?????00000??????????_??????,

    JR      = 32'b000000_????????????????????_001000,
    JALR    = 32'b000000_?????00000??????????_001001,
    J       = 32'b000010_????????????????????_??????,
    JAL     = 32'b000011_????????????????????_??????,

    LB      = 32'b100000_????????????????????_??????,
    LBU     = 32'b100100_????????????????????_??????,
    LH      = 32'b100001_????????????????????_??????,
    LHU     = 32'b100101_????????????????????_??????,
    LW      = 32'b100011_????????????????????_??????,
    SB      = 32'b101000_????????????????????_??????,
    SH      = 32'b101001_????????????????????_??????,
    SW      = 32'b101011_????????????????????_??????
} instruction_code_t;
`endif